module sd_reader(
	input					rst_n,
	input					clk,
	
	output		[7:0]		o_mm_data,
	output					o_mm_vld
);

endmodule

