// Code your design here
module draw_line(
  input					clk,
  
  input signed [15:0]	i_x1,
  input signed [15:0]	i_y1,
  input signed [15:0]	i_x2,
  input signed [15:0]	i_y2,
  
  output				rdy
);
  assign rdy = draw_state == DS_IDLE ? 1'b1 : 1'b0;
    
  reg signed [15:0] dx;
  reg signed [15:0] dy;
  
  assign dx = (i_x1 < i_x2) ? i_x2 - i_x1 : i_x1 - i_x2;
  assign dy = (i_y1 < i_y2) ? i_y2 - i_y1 : i_y1 - i_y2;
  
  wire swap_xy;
  assign swap_xy = (dx < dy) ? 1'b1 : 1'b0;
  
  reg signed [15:0] x1;
  reg signed [15:0] y1;
  reg signed [15:0] x2;
  reg signed [15:0] y2;
  
  assign x1 = swap_xy ? ((i_y1 < i_y2) ? i_y1 : i_y2) : ((i_x1 < i_x2) ? i_x1 : i_x2);
  assign x2 = swap_xy ? ((i_y1 < i_y2) ? i_y2 : i_y1) : ((i_x1 < i_x2) ? i_x2 : i_x1);
  assign y1 = swap_xy ? i_x1 : i_y1;
  assign y2 = swap_xy ? i_x2 : i_y2;
    
  reg signed [15:0] x;
  reg signed [15:0] y;
  reg signed [31:0] err;
  
  parameter [3:0] DS_NONE = 4'd0;
  parameter [3:0] DS_START = 4'd1;
  parameter [3:0] DS_DRAW = 4'd2;
  parameter [3:0] DS_IDLE = 4'd3;
  parameter [3:0] DS_STOP = 4'd4;
  
  reg [3:0] draw_state;
  
  initial draw_state = DS_NONE;
  
  always @ (posedge clk) begin
    case(draw_state)
      DS_NONE: begin
        $display("ds_none");
        draw_state <= DS_START;
      end
      DS_START: begin
        $display("ds_start dx=%d dy=%d", dx, dy);
        draw_state <= DS_DRAW;
        err <= -(dx / 2);
        x <= x1;
        y <= y1;
      end
      DS_DRAW: begin
        if(x <= x2) begin
          x <= x + 1;
          
          if(swap_xy) begin
            $display("swp put pixel (%d, %d)", y, x);
            
            err = err + dx;
            
            if(err >= 0) begin
              err <= err - dy;
              if(y1 < y2)
                y <= y + 1;
              else
                y <= y - 1;
            end
              
          end
          else begin
            $display("put pixel (%d, %d)", x, y);
          
            if(err + dy >= 0) begin
              err <= err + dy - dx;
              if(y1 < y2)
                y <= y + 1;
              else
                y <= y - 1;
            end
            else
              err <= err + dy;
          end
        end
        else begin
          draw_state <= DS_IDLE;
        end
      end
      DS_IDLE: begin
        draw_state <= DS_STOP;
        $display("idle state");
        //$finish;
      end      
    endcase
  end
  
endmodule

